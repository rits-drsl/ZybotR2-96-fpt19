/*
 MIT License

 Copyright (c) 2019 Yuya Kudo

 Permission is hereby granted, free of charge, to any person obtaining a copy
 of this software and associated documentation files (the "Software"), to deal
 in the Software without restriction, including without limitation the rights
 to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 copies of the Software, and to permit persons to whom the Software is
 furnished to do so, subject to the following conditions:

 The above copyright notice and this permission notice shall be included in all
 copies or substantial portions of the Software.

 THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 SOFTWARE.
 */

module general_cnt
  #(parameter
    INTERVAL = 100,
    localparam
    LB_INTERVAL = $clog2(INTERVAL))
   (output logic flag,
    input logic  clk,
    input logic  rstn);

   logic [LB_INTERVAL-1:0] cnt;

   always_comb begin
      flag = (cnt == INTERVAL - 1) ? 1 : 0;
   end

   always_ff @(posedge clk) begin
      if(rstn == 0) begin
         cnt <= 0;
      end
      else begin
         cnt <= cnt + 1;
         if(cnt == INTERVAL - 1) begin
            cnt <= 0;
         end
      end
   end
endmodule
